library verilog;
use verilog.vl_types.all;
entity t_scc_rom_mapper is
end t_scc_rom_mapper;
