library verilog;
use verilog.vl_types.all;
entity t_ch376 is
end t_ch376;
